present_val_reg: DFFSR PORT MAP(D=>n30, CLK=>clk, R=>n33, S=>1, Q=>stop_bit);
U2: OAI22X1 PORT MAP(A=>n28, B=>n32, C=>n3, D=>n31, Y=>n15);
Error: Bad Line.
U5: OAI22X1 PORT MAP(A=>n32, B=>n8, C=>n1, D=>n9, Y=>n19);
Error: Bad Line.
U9: OAI22X1 PORT MAP(A=>n32, B=>n6, C=>n1, D=>n7, Y=>n23);
Error: Bad Line.
U13: OAI22X1 PORT MAP(A=>n32, B=>n4, C=>n3, D=>n5, Y=>n27);
Error: Bad Line.
U17: NAND2X1 PORT MAP(A=>serial_in, B=>n3, Y=>n10);
Error: Bad Line.
U20: NAND2X1 PORT MAP(A=>packet_data0, B=>n32, Y=>n11);
Error: Bad Line.
U6: INVX4 PORT MAP(A=>n2, Y=>n1);
U8: INVX4 PORT MAP(A=>n2, Y=>n3);
U10: INVX8 PORT MAP(A=>shift_strobe, Y=>n32);
U12: INVX2 PORT MAP(A=>stop_bit, Y=>n4);
U14: INVX2 PORT MAP(A=>packet_data0, Y=>n5);
U15: INVX2 PORT MAP(A=>packet_data6, Y=>n6);
U18: INVX2 PORT MAP(A=>packet_data5, Y=>n7);
U21: INVX2 PORT MAP(A=>packet_data4, Y=>n8);
U22: INVX2 PORT MAP(A=>packet_data3, Y=>n9);
U32: INVX2 PORT MAP(A=>packet_data2, Y=>n28);
U33: INVX2 PORT MAP(A=>packet_data1, Y=>n31);
U34: INVX2 PORT MAP(A=>rst, Y=>n33);